module bram_ram_64 (
	input [15:0] in,
	input [5:0] address,
	input clk,
	input load,
	output [15:0] out
);

wire lda;
wire ldb;
wire ldc;
wire ldd;
wire lde;
wire ldf;
wire ldg;
wire ldh;
wire [15:0] outa;
wire [15:0] outb;
wire [15:0] outc;
wire [15:0] outd;
wire [15:0] oute;
wire [15:0] outf;
wire [15:0] outg;
wire [15:0] outh;

dmux_8_way dmux_8_way_a (
	.in(load),
	.select(address[5:3]),
	.a(lda),
	.b(ldb),
	.c(ldc),
	.d(ldd),
	.e(lde),
	.f(ldf),
	.g(ldg),
	.h(ldh)
);

bram_ram_8 bram_ram_8_a (
	.address(address[2:0]),
	.in(in),
	.clk(clk),
	.load(lda),
	.out(outa)
);
bram_ram_8 bram_ram_8_b (
	.address(address[2:0]),
	.in(in),
	.clk(clk),
	.load(ldb),
	.out(outb)
);
bram_ram_8 bram_ram_8_c (
	.address(address[2:0]),
	.in(in),
	.clk(clk),
	.load(ldc),
	.out(outc)
);
bram_ram_8 bram_ram_8_d (
	.address(address[2:0]),
	.in(in),
	.clk(clk),
	.load(ldd),
	.out(outd)
);
bram_ram_8 bram_ram_8_e (
	.in(in),
	.clk(clk),
	.load(lde),
	.out(oute)
);
bram_ram_8 bram_ram_8_f (
	.address(address[2:0]),
	.in(in),
	.clk(clk),
	.load(ldf),
	.out(outf)
);
bram_ram_8 bram_ram_8_g (
	.address(address[2:0]),
	.in(in),
	.clk(clk),
	.load(ldg),
	.out(outg)
);
bram_ram_8 bram_ram_8_h (
	.address(address[2:0]),
	.in(in),
	.clk(clk),
	.load(ldh),
	.out(outh)
);


n8WayMux16 n8WayMux16_a (
	.a(outa),
	.b(outb),
	.c(outc),
	.d(outd),
	.e(oute),
	.f(outf),
	.g(outg),
	.h(outh),
	.sel(address[5:3]),
	.out(out)
);



endmodule