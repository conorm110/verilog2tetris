module bram_ram_8 (
	input [15:0] in,
	input [2:0] address,
	input clk,
	input load,
	output [15:0] out
);



endmodule