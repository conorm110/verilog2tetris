module rzfpga_pc (

);



endmodule